`timescale 1ns / 1ps
module multu_tb;
	reg clk = 0;
	reg reset = 0;
	reg [31 : 0] a, b;
	wire [63 : 0] c;
	wire [63 : 0] rc;

	MULTU uut(.clk(clk), .reset(reset), .a(a), .b(b), .z(c));
    assign rc = a * b;

	always #5 clk = ~clk;
	initial begin
		reset <= 'b1;
		a <= 'b0;
		b <= 'b0;
		#5 reset <= 'b0;
		#30 a <= 'b0;
		b <= 'b11111111111111111111111111111111;
		#30 a <= 'b11111111111111111111111111111111;
		b <= 'b0;
		#30 a <= 'b11111111111111111111111111111111;
		b <= 'b11111111111111111111111111111111;
		#30 a <= 'b10000000000000000000000000000000;
		b <= 'b10101010101010101010101010101010;
		#30 a <= 'b10101010101010101010101010101010;
		b <= 'b10000000000000000000000000000000;
		#30 a <= 'b101101;
		b <= 'b1101000;
		#30 a <= 'b1000111;
		b <= 'b1110;
	end
endmodule
