`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/06/09 21:14:46
// Design Name: 
// Module Name: instr_dec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//指令译码器
module instr_dec(
    input [31 : 0] instr_code,
	output reg [31 : 0] instr_index
    );
	wire [11 : 0] temp;
	assign temp = {instr_code[31 : 26], instr_code[5 : 0]};
	always @ (*) begin
	    casez(temp)
		    //R-type
		    12'b000000100000: instr_index = 32'b00000000000000000000000000000001;//add
			12'b000000100001: instr_index = 32'b00000000000000000000000000000010;//addu
			12'b000000100010: instr_index = 32'b00000000000000000000000000000100;//sub
			12'b000000100011: instr_index = 32'b00000000000000000000000000001000;//subu
			12'b000000100100: instr_index = 32'b00000000000000000000000000010000;//and
			12'b000000100101: instr_index = 32'b00000000000000000000000000100000;//or
			12'b000000100110: instr_index = 32'b00000000000000000000000001000000;//xor
			12'b000000100111: instr_index = 32'b00000000000000000000000010000000;//nor
			12'b000000101010: instr_index = 32'b00000000000000000000000100000000;//slt
			12'b000000101011: instr_index = 32'b00000000000000000000001000000000;//sltu
			12'b000000000000: instr_index = 32'b00000000000000000000010000000000;//sll
			12'b000000000010: instr_index = 32'b00000000000000000000100000000000;//srl
			12'b000000000011: instr_index = 32'b00000000000000000001000000000000;//sra
			12'b000000000100: instr_index = 32'b00000000000000000010000000000000;//sllv
			12'b000000000110: instr_index = 32'b00000000000000000100000000000000;//srlv
			12'b000000000111: instr_index = 32'b00000000000000001000000000000000;//srav
			12'b000000001000: instr_index = 32'b00000000000000010000000000000000;//jr
			//I-type
			12'b001000??????: instr_index = 32'b00000000000000100000000000000000;//addi
			12'b001001??????: instr_index = 32'b00000000000001000000000000000000;//addiu
			12'b001100??????: instr_index = 32'b00000000000010000000000000000000;//andi
			12'b001101??????: instr_index = 32'b00000000000100000000000000000000;//ori
			12'b001110??????: instr_index = 32'b00000000001000000000000000000000;//xori
			12'b100011??????: instr_index = 32'b00000000010000000000000000000000;//lw
			12'b101011??????: instr_index = 32'b00000000100000000000000000000000;//sw
			12'b000100??????: instr_index = 32'b00000001000000000000000000000000;//beq
			12'b000101??????: instr_index = 32'b00000010000000000000000000000000;//bne
			12'b001010??????: instr_index = 32'b00000100000000000000000000000000;//slti
			12'b001011??????: instr_index = 32'b00001000000000000000000000000000;//sltiu
			12'b001111??????: instr_index = 32'b00010000000000000000000000000000;//lui
			//J-type
			12'b000010??????: instr_index = 32'b00100000000000000000000000000000;//j
			12'b000011??????: instr_index = 32'b01000000000000000000000000000000;//jal
			default:          instr_index = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
		endcase
	end			
endmodule
